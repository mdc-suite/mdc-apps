`ifndef LAYERS_SIZES_VH
`define LAYERS_SIZES_VH
	`define kern_s_0	16*3*1
	`define kern_s_k_0	16
	`define kern_s_1	16*3*1
	`define kern_s_k_1	16
	`define kern_s_2	8*3*1
	`define kern_s_k_2	8
	`define kern_s_3	16*8*9
	`define kern_s_k_3	16
	`define kern_s_4	8*3*1
	`define kern_s_k_4	8
	`define kern_s_5	16*8*9
	`define kern_s_k_5	16
	`define kern_s_6	16*16*9
	`define kern_s_k_6	16
	`define kern_s_7	32*64*1	
	`define kern_s_k_7	32
	`define kern_s_8	32*64*1	
	`define kern_s_k_8	32
	`define kern_s_9	16*64*1	
	`define kern_s_k_9	16
	`define kern_s_10	32*16*9	
	`define kern_s_k_10	32
	`define kern_s_11	16*64*1	
	`define kern_s_k_11	16
	`define kern_s_12	32*16*9
	`define kern_s_k_12	32
	`define kern_s_13	32*32*9	
	`define kern_s_k_13	32
	`define kern_s_14	64*128*1	
	`define kern_s_k_14	64
	`define kern_s_15	64*128*1	
	`define kern_s_k_15	64
	`define kern_s_16	32*128*1	
	`define kern_s_k_16	32
	`define kern_s_17	64*32*9	
	`define kern_s_k_17	64
	`define kern_s_18	32*128*1	
	`define kern_s_k_18	32
	`define kern_s_19	64*32*9		
	`define kern_s_k_19	64
	`define kern_s_20	64*64*9		
	`define kern_s_k_20	64
	`define kern_s_21	16*256*1	
	`define kern_s_k_21	16
`endif