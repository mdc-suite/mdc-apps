`ifndef MY_TYPES_VH
`define MY_TYPES_VH
	`define data_width 16
	`define coeff_width 8
`endif